// MIT License

// Copyright (c) 2020 Jonghoon Won (jonghoon@gatech.edu)

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.


import Fifo::*;


typedef Bit#(64) Data;


interface Adder;
    method Action putA(Data data);
    method Action putB(Data data);
    method ActionValue#(Data) getResult();
endinterface


(* synthesize *)
module mkAdder(Adder);
    Fifo#(1, Data) argA <- mkPipelineFifo;
    Fifo#(1, Data) argB <- mkPipelineFifo;
    Fifo#(1, Data) result <- mkBypassFifo;


    rule doAddition;
        let a = argA.first;
        let b = argB.first;
        argA.deq;
        argB.deq;

        result.enq(a + b);
    endrule


    method Action putA(Data data);
        argA.enq(data);
    endmethod

    method Action putB(Data data);
        argB.enq(data);
    endmethod

    method ActionValue#(Data) getResult();
        result.deq;
        return result.first;
    endmethod
endmodule
